module Top_Module (
    input clk,
    input reset,
    input [15:0] soil_voltage_mv,
    input [15:0] dht11_voltage_mv,
    input [15:0] rain_voltage_mv,
    input [3:0] keypad_row,
    input [3:0] keypad_col,
    output keypad_start,
    output keypad_accept,
    output keypad_backspace,
    output [3:0] category,
    output [9:0] new_value,
    output pump_on,
    output rain_present,
    output watering_in_progress,
    output sensor_enable,
    output sda,
    output scl,
    output [9:0] soil_digital,
    output [9:0] dht11_digital,
    output [9:0] rain_digital,
    output [7:0] irrigation_time,
    output [9:0] new_soil_dry,
    output [9:0] new_soil_moist,
    output [9:0] new_soil_wet,
    output [9:0] new_temp_cold,
    output [9:0] new_temp_warm,
    output [9:0] new_temp_hot,
    output [9:0] new_rain_no,
    output [9:0] new_rain_yes,
    output update_soil_dry,
    output update_soil_moist,
    output update_soil_wet,
    output update_temp_cold,
    output update_temp_warm,
    output update_temp_hot,
    output update_rain_no,
    output update_rain_yes,
    output updated,
    output [7:0] watering_timer,
    output [9:0] param_soil_dry,
    output [9:0] param_soil_moist,
    output [9:0] param_soil_wet,
    output [9:0] param_temp_cold,
    output [9:0] param_temp_warm,
    output [9:0] param_temp_hot,
    output [9:0] param_rain_no,
    output [9:0] param_rain_yes,
    output [23:0] lcd_data,
    output [23:0] lcd_message_data
);

    ADC_SENSOR uut_adc (
        .clk(clk),
        .reset(reset),
        .soil_voltage_mv(soil_voltage_mv),
        .dht11_voltage_mv(dht11_voltage_mv),
        .rain_voltage_mv(rain_voltage_mv),
        .sensor_enable(sensor_enable),
        .soil_digital(soil_digital),
        .dht11_digital(dht11_digital),
        .rain_digital(rain_digital)
    );

    FUZZIFIKASI uut_fuzzy (
        .clk(clk),
        .reset(reset),
        .new_soil_dry(new_soil_dry),
        .new_soil_moist(new_soil_moist),
        .new_soil_wet(new_soil_wet),
        .new_temp_cold(new_temp_cold),
        .new_temp_warm(new_temp_warm),
        .new_temp_hot(new_temp_hot),
        .new_rain_no(new_rain_no),
        .new_rain_yes(new_rain_yes),
        .update_soil_dry(update_soil_dry),
        .update_soil_moist(update_soil_moist),
        .update_soil_wet(update_soil_wet),
        .update_temp_cold(update_temp_cold),
        .update_temp_warm(update_temp_warm),
        .update_temp_hot(update_temp_hot),
        .update_rain_no(update_rain_no),
        .update_rain_yes(update_rain_yes),
        .soil_digital(soil_digital),
        .dht11_digital(dht11_digital),
        .rain_digital(rain_digital),
        .irrigation_time(irrigation_time),
        .rain_present(rain_present),
        .PARAM_SOIL_DRY(param_soil_dry),
        .PARAM_SOIL_MOIST(param_soil_moist),
        .PARAM_SOIL_WET(param_soil_wet),
        .PARAM_TEMP_COLD(param_temp_cold),
        .PARAM_TEMP_WARM(param_temp_warm),
        .PARAM_TEMP_HOT(param_temp_hot),
        .PARAM_RAIN_NO(param_rain_no),
        .PARAM_RAIN_YES(param_rain_yes)
    );

    Penyiraman_Otomatis uut_pump (
        .clk(clk),
        .reset(reset),
        .irrigation_time(irrigation_time),
        .pump_on(pump_on),
        .sensor_enable(sensor_enable),
        .watering_in_progress(watering_in_progress),
        .watering_timer(watering_timer)
    );


    KEYPAD4x4 uut_keypad (
        .clk(clk),
        .reset(reset),
        .keypad_row(keypad_row),
        .keypad_col(keypad_col),
		  .category(category),
		  .new_value(new_value),
        .start(keypad_start),
        .accept(keypad_accept),
        .backspace(keypad_backspace),
        .PARAM_SOIL_DRY(param_soil_dry),
        .PARAM_SOIL_MOIST(param_soil_moist),
        .PARAM_SOIL_WET(param_soil_wet),
        .PARAM_TEMP_COLD(param_temp_cold),
        .PARAM_TEMP_WARM(param_temp_warm),
        .PARAM_TEMP_HOT(param_temp_hot),
        .PARAM_RAIN_NO(param_rain_no),
        .PARAM_RAIN_YES(param_rain_yes),
        .updated(updated),
        .NEW_PARAM_SOIL_DRY(new_soil_dry),
        .NEW_PARAM_SOIL_MOIST(new_soil_moist),
        .NEW_PARAM_SOIL_WET(new_soil_wet),
        .NEW_PARAM_TEMP_COLD(new_temp_cold),
        .NEW_PARAM_TEMP_WARM(new_temp_warm),
        .NEW_PARAM_TEMP_HOT(new_temp_hot),
        .NEW_PARAM_RAIN_NO(new_rain_no),
        .NEW_PARAM_RAIN_YES(new_rain_yes),
        .update_soil_dry(update_soil_dry),
        .update_soil_moist(update_soil_moist),
        .update_soil_wet(update_soil_wet),
        .update_temp_cold(update_temp_cold),
        .update_temp_warm(update_temp_warm),
        .update_temp_hot(update_temp_hot),
        .update_rain_no(update_rain_no),
        .update_rain_yes(update_rain_yes)
    );

    LCD_I2C uut_lcd (
        .clk(clk),
        .reset(reset),
        .dht11_digital(dht11_digital),
        .soil_digital(soil_digital),
        .rain_digital(rain_digital),
        .watering_in_progress(watering_in_progress),
        .watering_timer(watering_timer),
        .sensor_enable(sensor_enable),
        .lcd_data(lcd_data),
        .lcd_message_data(lcd_message_data),
        .sda(sda),
        .scl(scl)
    );

endmodule
